package ring_pkg;

    import uvm_pkg::*;

`include "uvm_macros.svh"

`include "ring_transaction.sv"


`include "ring_monitor.sv"
`include "ring_sequencer.sv"
`include "ring_driver.sv"
`include "ring_agent.sv"
`include "ring_sequence.sv"




endpackage
