package hello_pkg;

    import uvm_pkg::*;

`include "uvm_macros.svh"

`include "hello_transaction.sv"


`include "hello_monitor.sv"
`include "hello_sequencer.sv"
`include "hello_driver.sv"
`include "hello_agent.sv"
`include "hello_sequence.sv"




endpackage
